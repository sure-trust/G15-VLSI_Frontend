display from top
display from test
display from environment
display from generator
d_in=11011100,done=0,ss=0,mosi=0
display from driver
d_in=11011100,done=0,ss=0,mosi=0
display from monitor
d_in=11011100,done=0,ss=0,mosi=0
scoreboard
matched outputs
state=0
state=0
display from monitor
d_in=11011100,done=0,ss=1,mosi=0
scoreboard
matched outputs
state=0
state=0
display from monitor
d_in=11011100,done=0,ss=1,mosi=0
scoreboard
matched outputs
state=0
state=0
display from monitor
d_in=11011100,done=0,ss=1,mosi=0
scoreboard
matched outputs
state=0
state=0
display from monitor
d_in=11011100,done=0,ss=1,mosi=0
scoreboard
matched outputs
state=0
state=0
$finish called from file "testbench.sv", line 30.
$finish at simulation time                   20
           V C S   S i m u l a t i o n   R e p o r t 
Time: 20 ns
CPU Time:      0.640 seconds;       Data structure size:   0.0Mb
Tue Mar 19 23:52:14 2024
Finding VCD file...
./dump.vcd