//Counter
module counter(clk1,rst1,A,clk2,rst2,B);
  input clk1,clk2,rst1,rst2;
  output reg [3:0]A,B;
  
  counterA dut1(clk1,rst1,A);
  
  and a1(clk2,A[0],A[1]);
  
  counterB dut2(clk2,rst2,B);
  
endmodule

//counter A

module counterA (
  input wire clk,
  input wire reset,
  output reg [3:0] count
);

  always @(posedge clk or posedge reset) begin
    if (reset)
      count <= 4'b0000;
    else
      count <= count + 1;
  end

endmodule

//counter B

module CounterB (
  input wire clk,
  input wire reset,
  output reg [3:0] count
);

  always @(posedge clk or posedge reset) begin
    if (reset)
      count <= 4'b1111;
    else
      count <= count - 1;
  end

endmodule


//test bench

module tb_counter;

  reg clk1, rst1, clk2, rst2;
  wire [3:0] A, B;

  
  counter dut(
    .clk1(clk1),
    .rst1(rst1),
    .A(A),
    .clk2(clk2),
    .rst2(rst2),
    .B(B)
  );

  
  initial begin
    clk1 = 0;
    forever #5 clk1 = ~clk1; 
  end

  initial begin
    clk2 = 0;
    forever #10 clk2 = ~clk2;  
  end

 
  initial begin
    rst1 = 1; rst2 = 1; 
    #15 rst1 = 0; rst2 = 0;   units

    
    $monitor("Time=%0t: A=%b, B=%b", $time, A, B);

   
    #100 $finish;
  end

endmodule

