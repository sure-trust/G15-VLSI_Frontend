`include "uvm_macros.svh"
import uvm_pkg::*;
`include "interface.sv"
`include "sequence_item.sv"
`include "sequence1.sv"
`include "sequence2.sv"
`include "sequence3.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "agent.sv"
`include "environment.sv"
`include "test.sv"