interface intf(input logic clk,rst);
  
  logic [1:0] addr;
  logic wr_en;
  logic rd_en;
  logic [7:0] wdata;
  logic [7:0] rdata;
   clocking driv_cb@(posedge clk);
  default input #1 output #2;
    output addr;
     output wr_en;
     output rd_en;
     output wdata;
    input rdata;
    
  endclocking
  
  clocking mon_cb@(posedge clk);
    input addr;
    input wr_en;
    input rd_en;
    input wdata;
    input rdata;
  endclocking
  
  endinterface