`include "uvm_macros.svh"
 import uvm_pkg::*;

`include "interface.sv"
`include "sequence_item.sv"
`include "sequence.sv"
//`include "sequnecer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "environment.sv"
`include "test.sv"
/////////////build the seq for random length with and without priority

////////////////////////////////////////////////////////////////////////////////////
