// Design code
module seq_detector_1010(input bit clk, rst_n, x, output z);
  parameter A = 4'h1;
  parameter B = 4'h2;
  parameter C = 4'h3;
  parameter D = 4'h4;
  
  bit [3:0] state, next_state;
  always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin 
      state <= A;
    end
    else state <= next_state;
  end
  
  always @(state or x) begin
    case(state)
      A: begin
        if(x == 0) next_state = B;
           else       next_state = A;
         end
      B: begin
        if(x == 1) next_state = C;
           else       next_state = B;
         end
      C: begin
        if(x == 1) next_state = D;
           else       next_state = B;
         end
      D: begin
        if(x == 0) next_state = A; 
           else       next_state = A;
         end
      default: next_state = A;
    endcase
  end
  assign z = (state == D) && (x == 0)? 1:0;
endmodule


//Test Bench

module TB;
  reg clk, rst_n, x;
  wire z;
  
  seq_detector_1010 sd(clk, rst_n, x, z);
  initial clk = 0;   
  always #2 clk = ~clk;
    
  initial begin
    x = 0;
    #1 rst_n = 0;
    #2 rst_n = 1;
     #4 x = 0;
    #4 x = 1;
    #4 x = 1;
    #4 x = 1;
    
    #4 x = 0;
    #4 x = 1;
    #4 x = 1;
    #4 x = 0;
    
   
  
    #10;
    $finish;
  end
  
  initial begin
    // Dump waves
    $dumpfile("dump.vcd");
    $dumpvars(0);
  end
endmodule
